`ifndef _{:UPPERNAME:}_SEQUENCER_SV_
`define _{:UPPERNAME:}_SEQUENCER_SV_

typedef uvm_sequencer #({:NAME:}_seq_item) {:NAME:}_sequencer;

`endif

